parameter WORD_SIZE = 16;

`define ALU_ADD 4'h0 //0000
`define ALU_SUB 4'h1
`define ALU_MUL 4'h2
`define ALU_SLT 4'h3
`define ALU_AND 4'h4
`define ALU_OR 4'h5
`define ALU_XOR 4'h6
`define ALU_SHL 4'h7 
`define ALU_SHR 4'h8 //1000