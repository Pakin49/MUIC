parameter WORD_SIZE = 16;

`define ALU_ADD 3'h0 //000
`define ALU_SUB 3'h1
`define ALU_MUL 3'h2
`define ALU_SLT 3'h3
`define ALU_AND 3'h4
`define ALU_OR 3'h5
`define ALU_XOR 3'h6
`define ALU_SHIFT 3'h7 //111